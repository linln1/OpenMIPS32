module  id(

    input wire              rst,
    input wire['InstAddrBus]              pc_i,
    input wire['InstBus]                  inst_i,
    
    // 读取的Regfile的值
    input wire['RegBus]                   reg1_data_i,
    input wire['RegBus]                   reg2_data_i,
    
    // 输出的Regfile的值 
    output reg                            reg1_read_o,
    output reg                            reg2_read_o,
    
    output reg['RegAddrBus]               reg1_addr_o,
    output reg['RegAddrBus]               reg2_addr_o,
    
    // 送到执行阶段的信息
    output reg['AluOpBus]                 aluop_o,
    output reg['AluSelBus]                 alusel_o,
    output reg['RegBus]                 reg1_o,
    output reg['RegBus]                 reg2_o,
    output reg['RegAddrBus]                 wd_o,
    output reg                            wreg_o,
);


//取得指令的指令码，功能码
//对于ori指令只需要通过判断26-31bit的值，即可判断是否ori指令
wire[5:0]   op  =   inst_i[31:26];
wire[4:0]   op2 =   inst_i[10:6];
wire[5:0]   op3 =   inst_i[5:0];
wire[4:0]   op4 =   inst_i[20:16];
//保存指令执行需要的立即数
reg['RegBus]    imm;
//指示指令是否有效
reg instvalid;


/***************************************************
                第一段:译码
****************************************************/
    always  @   (*) begin
        if  (rst == 'RstEnable) begin
            aluop_o     <=      'EXE_NOP_OP;
            alusel_o    <=      'EXE_RES_NOP;
            wd_o        <=      'NOPRegAddr;
            wreg_o      <=      'WriteDisable;
            instvalid   <=      'InstValid;
            reg1_read_o <=      1'b0;
            reg2_read_o <=      1'b0;
            reg1_addr_o <=      'NOPRegAddr;
            reg2_addr_o <=      'NOPRegAddr;
            imm         <=      32'h0;
        end else    begin
            aluop_o     <=      'EXE_NOP_OP;
            alusel_o    <=      'EXE_RES_NOP;
            wd_o        <=      inst_i[15:11];
            wreg_o      <=      'WriteDisable;
            instvalid   <=      'InstValid;
            reg1_read_o <=      1'b0;
            reg2_read_o <=      1'b0;
            reg1_addr_o <=      'inst_i[25:21];
            reg2_addr_o <=      'inst_i[20:16];
            imm         <=      'ZeroWord;


            case(op):
                'EXE_ORI:       begin
                    wreg_o      <=      'WriteEnable;
                    aluop_o     <=      'EXE_OR_OP;
                    alusel_o    <=      'EXE_RES_LOGIC;
                    reg1_read_o <=      1'b1;
                    reg2_read_o <=      1'b0;
                    imm         <=      {16'h0, inst_i[15:0]}
                    wd_o        <=      inst_i[20:16];
                    instvalid   <=      'InstValid;
                end
                
                default:begin
                end
                end
            endcase
            
        end
    end
      
/***************************************************
                第2段:确定运算的源操作数1
****************************************************/
    always  @   (*)     begin
        if  (rst ==  'RstEnable)    begin
                reg1_o  <=  'ZeroWord;
        end else if (reg1_read_o  ==  1'b1) begin
                reg1_o <=  reg1_data_i;
        end else if (reg1_read_o  ==  1'b0) begin
                reg1_o <=  imm;
        end else begin
                reg1_o <= 'ZeroWord;
        end
    end
/***************************************************
                第3段:确定运算的源操作数2
****************************************************/
    always  @   (*)     begin
        if  (rst == 'RstEnable)     begin
                reg2_o  <=  'ZeroWord;
        end else if (reg2_read_o == 1'b1) begin
                reg2_o  <=  reg2_data_i;
        end else if (reg2_read_o == 1'b0) begin
                reg2_o  <=  imm;
        end else begin
                reg2_o  <=  'ZeroWord;
        end
    end
    
endmodule


